module crud