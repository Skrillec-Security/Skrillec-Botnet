module server