module attack_system


pub fn send_attack(ip string, port string, time string, method string) int {

}

pub fn fill_api(ip string, port string, time string, method string) {

}

pub fn get_all_api() {
	
}