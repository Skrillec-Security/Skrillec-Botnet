module server

pub fn bot_attack() { 
	
}