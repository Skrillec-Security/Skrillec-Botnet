module skrillec_cp

import os

pub fn main_cp() {
	for {
		mut input_cmd := os.input(">>> ")
		
	}
}