module server

import net
import net.http

pub fn validate_token(token string) {

}