module attack_system


pub fn send_attack(ip string, port string, time string, method string) {
	
}