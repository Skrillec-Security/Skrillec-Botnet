module crud

import mysql

// pub fn total_users(mut s mysql.Connection) int {
	
// }