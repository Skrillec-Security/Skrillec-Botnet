module config

pub struct AppInfo{
	pub mut:
		title		string = "Skrillec Botnet"
		description	string = "The New 2022 All-In-One Botnet. Eliminating the hassle of looking for all botnet related files to start one up!"
		version		string = "4.00"
}