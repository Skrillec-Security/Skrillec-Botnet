module attack_system
