module crud

import crud
import mysql

pub fn get_user(username string, mut s mysql.Connection) {
	rows := crud.get_row()
}