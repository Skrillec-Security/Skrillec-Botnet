module config

pub fn get_net_info() []string {

}