module utils