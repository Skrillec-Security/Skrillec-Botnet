module utils

