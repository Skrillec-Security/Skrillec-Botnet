module crud

