module config

pub struct AppInfo{
	pub mut:
		title		string = "Skrillec Botnet"
		description	string = "The New 2022 All-In-One Botnet. Eliminating the hassle of looking for all botnet related files to start one up!"
		version		string = "4.00"
}

const (
	//Colors
	Default			= ""
	Black			= ""
	Red				= ""
	Green			= ""
	Yellow			= ""
	Blue			= ""
	Purple			= ""
	Cyan			= ""
	Light_Grey		= ""
	Dark_Grey		= ""
	Light_red		= ""
	Light_Green		= ""
	Light_Yellow	= ""
	Light_Blue		= ""
	Light_Purple	= ""
	Light_Cyan		= ""
	White			= ""
	// Background Colors
	Default_BG		= ""
	Black_BG		= ""
	Red_BG			= ""
	Green_BG		= ""
	Yellow_BG		= ""
	Blue_BG			= ""
	Purple_BG		= ""
	Cyan_BG			= ""
)